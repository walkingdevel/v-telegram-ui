module users

pub struct User {
pub:
	username    string
	fullname    string
	avatar_path string
}
